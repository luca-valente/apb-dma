`define NUM_REGS 6
